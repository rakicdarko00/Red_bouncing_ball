library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Tue May 16 17:29:36 2017

	signal mem : ram_t := (


--			***** 8x8 IMAGES *****

--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"001859DE", -- R: 222 G: 89 B: 24
		2 =>	x"00E2F2FF", -- R: 255 G: 242 B: 226
		3 =>	x"00EAD999", -- R: 153 G: 217 B: 234
		4 =>	x"00429DFB", -- R: 251 G: 157 B: 66
		5 =>	x"003496FC", -- R: 252 G: 150 B: 52
		6 =>	x"003A9DFF", -- R: 255 G: 157 B: 58
		7 =>	x"003B9DFF", -- R: 255 G: 157 B: 59
		8 =>	x"003599FF", -- R: 255 G: 153 B: 53
		9 =>	x"004B91C0", -- R: 192 G: 145 B: 75
		10 =>	x"00947C00", -- R: 0 G: 124 B: 148
		11 =>	x"00877D00", -- R: 0 G: 125 B: 135
		12 =>	x"008E860E", -- R: 14 G: 134 B: 142
		13 =>	x"003B9AFC", -- R: 252 G: 154 B: 59
		14 =>	x"00399DFF", -- R: 255 G: 157 B: 57
		15 =>	x"001C68DB", -- R: 219 G: 104 B: 28
		16 =>	x"001E6CDE", -- R: 222 G: 108 B: 30
		17 =>	x"003495FF", -- R: 255 G: 149 B: 52
		18 =>	x"003F96E6", -- R: 230 G: 150 B: 63
		19 =>	x"005A8D8E", -- R: 142 G: 141 B: 90
		20 =>	x"007C821E", -- R: 30 G: 130 B: 124
		21 =>	x"008C8100", -- R: 0 G: 129 B: 140
		22 =>	x"00208BFB", -- R: 251 G: 139 B: 32
		23 =>	x"003697FC", -- R: 252 G: 151 B: 54
		24 =>	x"003CA0FF", -- R: 255 G: 160 B: 60
		25 =>	x"000540C0", -- R: 192 G: 64 B: 5
		26 =>	x"000846C4", -- R: 196 G: 70 B: 8
		27 =>	x"00043FC1", -- R: 193 G: 63 B: 4
		28 =>	x"003491F7", -- R: 247 G: 145 B: 52
		29 =>	x"003799FF", -- R: 255 G: 153 B: 55
		30 =>	x"002C9BFF", -- R: 255 G: 155 B: 44
		31 =>	x"00728640", -- R: 64 G: 134 B: 114
		32 =>	x"00897E00", -- R: 0 G: 126 B: 137
		33 =>	x"007A7000", -- R: 0 G: 112 B: 122
		34 =>	x"00218CFB", -- R: 251 G: 140 B: 33
		35 =>	x"002B91FB", -- R: 251 G: 145 B: 43
		36 =>	x"001C68DA", -- R: 218 G: 104 B: 28
		37 =>	x"000035B8", -- R: 184 G: 53 B: 0
		38 =>	x"0041A8FF", -- R: 255 G: 168 B: 65
		39 =>	x"003DA0FF", -- R: 255 G: 160 B: 61
		40 =>	x"0034A3FF", -- R: 255 G: 163 B: 52
		41 =>	x"008C8000", -- R: 0 G: 128 B: 140
		42 =>	x"007E831C", -- R: 28 G: 131 B: 126
		43 =>	x"00309AFF", -- R: 255 G: 154 B: 48
		44 =>	x"003399FF", -- R: 255 G: 153 B: 51
		45 =>	x"00577AB9", -- R: 185 G: 122 B: 87
		46 =>	x"00807700", -- R: 0 G: 119 B: 128
		47 =>	x"007A7100", -- R: 0 G: 113 B: 122
		48 =>	x"003898FC", -- R: 252 G: 152 B: 56
		49 =>	x"001F6DDE", -- R: 222 G: 109 B: 31
		50 =>	x"00043EBE", -- R: 190 G: 62 B: 4
		51 =>	x"002F9AFF", -- R: 255 G: 154 B: 47
		52 =>	x"00848109", -- R: 9 G: 129 B: 132
		53 =>	x"003698FF", -- R: 255 G: 152 B: 54
		54 =>	x"003B97EF", -- R: 239 G: 151 B: 59
		55 =>	x"0033A2FF", -- R: 255 G: 162 B: 51
		56 =>	x"00269DFF", -- R: 255 G: 157 B: 38
		57 =>	x"008A7F00", -- R: 0 G: 127 B: 138
		58 =>	x"002E9AFF", -- R: 255 G: 154 B: 46
		59 =>	x"008D7E00", -- R: 0 G: 126 B: 141
		60 =>	x"003F95E4", -- R: 228 G: 149 B: 63
		61 =>	x"003598FF", -- R: 255 G: 152 B: 53
		62 =>	x"003C9AFC", -- R: 252 G: 154 B: 60
		63 =>	x"003199FF", -- R: 255 G: 153 B: 49
		64 =>	x"0069885F", -- R: 95 G: 136 B: 105
		65 =>	x"00658A6C", -- R: 108 G: 138 B: 101
		66 =>	x"006A895E", -- R: 94 G: 137 B: 106
		67 =>	x"003997F7", -- R: 247 G: 151 B: 57
		68 =>	x"003E95E8", -- R: 232 G: 149 B: 62
		69 =>	x"003299FF", -- R: 255 G: 153 B: 50
		70 =>	x"003499FF", -- R: 255 G: 153 B: 52
		71 =>	x"004A91C0", -- R: 192 G: 145 B: 74
		72 =>	x"00E8A200", -- R: 0 G: 162 B: 232
		73 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		74 =>	x"00584000", -- R: 0 G: 64 B: 88
		75 =>	x"00C9DDFF", -- R: 255 G: 221 B: 201
		76 =>	x"000038F8", -- R: 248 G: 56 B: 0
		77 =>	x"00007CAC", -- R: 172 G: 124 B: 0
		78 =>	x"0040A4FF", -- R: 255 G: 164 B: 64
		79 =>	x"00349DEF", -- R: 239 G: 157 B: 52
		80 =>	x"003092E0", -- R: 224 G: 146 B: 48
		81 =>	x"00309AEA", -- R: 234 G: 154 B: 48
		82 =>	x"00000000", -- R: 0 G: 0 B: 0
		83 =>	x"00000000", -- R: 0 G: 0 B: 0
		84 =>	x"00000000", -- R: 0 G: 0 B: 0
		85 =>	x"00000000", -- R: 0 G: 0 B: 0
		86 =>	x"00000000", -- R: 0 G: 0 B: 0
		87 =>	x"00000000", -- R: 0 G: 0 B: 0
		88 =>	x"00000000", -- R: 0 G: 0 B: 0
		89 =>	x"00000000", -- R: 0 G: 0 B: 0
		90 =>	x"00000000", -- R: 0 G: 0 B: 0
		91 =>	x"00000000", -- R: 0 G: 0 B: 0
		92 =>	x"00000000", -- R: 0 G: 0 B: 0
		93 =>	x"00000000", -- R: 0 G: 0 B: 0
		94 =>	x"00000000", -- R: 0 G: 0 B: 0
		95 =>	x"00000000", -- R: 0 G: 0 B: 0
		96 =>	x"00000000", -- R: 0 G: 0 B: 0
		97 =>	x"00000000", -- R: 0 G: 0 B: 0
		98 =>	x"00000000", -- R: 0 G: 0 B: 0
		99 =>	x"00000000", -- R: 0 G: 0 B: 0
		100 =>	x"00000000", -- R: 0 G: 0 B: 0
		101 =>	x"00000000", -- R: 0 G: 0 B: 0
		102 =>	x"00000000", -- R: 0 G: 0 B: 0
		103 =>	x"00000000", -- R: 0 G: 0 B: 0
		104 =>	x"00000000", -- R: 0 G: 0 B: 0
		105 =>	x"00000000", -- R: 0 G: 0 B: 0
		106 =>	x"00000000", -- R: 0 G: 0 B: 0
		107 =>	x"00000000", -- R: 0 G: 0 B: 0
		108 =>	x"00000000", -- R: 0 G: 0 B: 0
		109 =>	x"00000000", -- R: 0 G: 0 B: 0
		110 =>	x"00000000", -- R: 0 G: 0 B: 0
		111 =>	x"00000000", -- R: 0 G: 0 B: 0
		112 =>	x"00000000", -- R: 0 G: 0 B: 0
		113 =>	x"00000000", -- R: 0 G: 0 B: 0
		114 =>	x"00000000", -- R: 0 G: 0 B: 0
		115 =>	x"00000000", -- R: 0 G: 0 B: 0
		116 =>	x"00000000", -- R: 0 G: 0 B: 0
		117 =>	x"00000000", -- R: 0 G: 0 B: 0
		118 =>	x"00000000", -- R: 0 G: 0 B: 0
		119 =>	x"00000000", -- R: 0 G: 0 B: 0
		120 =>	x"00000000", -- R: 0 G: 0 B: 0
		121 =>	x"00000000", -- R: 0 G: 0 B: 0
		122 =>	x"00000000", -- R: 0 G: 0 B: 0
		123 =>	x"00000000", -- R: 0 G: 0 B: 0
		124 =>	x"00000000", -- R: 0 G: 0 B: 0
		125 =>	x"00000000", -- R: 0 G: 0 B: 0
		126 =>	x"00000000", -- R: 0 G: 0 B: 0
		127 =>	x"00000000", -- R: 0 G: 0 B: 0
		128 =>	x"00000000", -- R: 0 G: 0 B: 0
		129 =>	x"00000000", -- R: 0 G: 0 B: 0
		130 =>	x"00000000", -- R: 0 G: 0 B: 0
		131 =>	x"00000000", -- R: 0 G: 0 B: 0
		132 =>	x"00000000", -- R: 0 G: 0 B: 0
		133 =>	x"00000000", -- R: 0 G: 0 B: 0
		134 =>	x"00000000", -- R: 0 G: 0 B: 0
		135 =>	x"00000000", -- R: 0 G: 0 B: 0
		136 =>	x"00000000", -- R: 0 G: 0 B: 0
		137 =>	x"00000000", -- R: 0 G: 0 B: 0
		138 =>	x"00000000", -- R: 0 G: 0 B: 0
		139 =>	x"00000000", -- R: 0 G: 0 B: 0
		140 =>	x"00000000", -- R: 0 G: 0 B: 0
		141 =>	x"00000000", -- R: 0 G: 0 B: 0
		142 =>	x"00000000", -- R: 0 G: 0 B: 0
		143 =>	x"00000000", -- R: 0 G: 0 B: 0
		144 =>	x"00000000", -- R: 0 G: 0 B: 0
		145 =>	x"00000000", -- R: 0 G: 0 B: 0
		146 =>	x"00000000", -- R: 0 G: 0 B: 0
		147 =>	x"00000000", -- R: 0 G: 0 B: 0
		148 =>	x"00000000", -- R: 0 G: 0 B: 0
		149 =>	x"00000000", -- R: 0 G: 0 B: 0
		150 =>	x"00000000", -- R: 0 G: 0 B: 0
		151 =>	x"00000000", -- R: 0 G: 0 B: 0
		152 =>	x"00000000", -- R: 0 G: 0 B: 0
		153 =>	x"00000000", -- R: 0 G: 0 B: 0
		154 =>	x"00000000", -- R: 0 G: 0 B: 0
		155 =>	x"00000000", -- R: 0 G: 0 B: 0
		156 =>	x"00000000", -- R: 0 G: 0 B: 0
		157 =>	x"00000000", -- R: 0 G: 0 B: 0
		158 =>	x"00000000", -- R: 0 G: 0 B: 0
		159 =>	x"00000000", -- R: 0 G: 0 B: 0
		160 =>	x"00000000", -- R: 0 G: 0 B: 0
		161 =>	x"00000000", -- R: 0 G: 0 B: 0
		162 =>	x"00000000", -- R: 0 G: 0 B: 0
		163 =>	x"00000000", -- R: 0 G: 0 B: 0
		164 =>	x"00000000", -- R: 0 G: 0 B: 0
		165 =>	x"00000000", -- R: 0 G: 0 B: 0
		166 =>	x"00000000", -- R: 0 G: 0 B: 0
		167 =>	x"00000000", -- R: 0 G: 0 B: 0
		168 =>	x"00000000", -- R: 0 G: 0 B: 0
		169 =>	x"00000000", -- R: 0 G: 0 B: 0
		170 =>	x"00000000", -- R: 0 G: 0 B: 0
		171 =>	x"00000000", -- R: 0 G: 0 B: 0
		172 =>	x"00000000", -- R: 0 G: 0 B: 0
		173 =>	x"00000000", -- R: 0 G: 0 B: 0
		174 =>	x"00000000", -- R: 0 G: 0 B: 0
		175 =>	x"00000000", -- R: 0 G: 0 B: 0
		176 =>	x"00000000", -- R: 0 G: 0 B: 0
		177 =>	x"00000000", -- R: 0 G: 0 B: 0
		178 =>	x"00000000", -- R: 0 G: 0 B: 0
		179 =>	x"00000000", -- R: 0 G: 0 B: 0
		180 =>	x"00000000", -- R: 0 G: 0 B: 0
		181 =>	x"00000000", -- R: 0 G: 0 B: 0
		182 =>	x"00000000", -- R: 0 G: 0 B: 0
		183 =>	x"00000000", -- R: 0 G: 0 B: 0
		184 =>	x"00000000", -- R: 0 G: 0 B: 0
		185 =>	x"00000000", -- R: 0 G: 0 B: 0
		186 =>	x"00000000", -- R: 0 G: 0 B: 0
		187 =>	x"00000000", -- R: 0 G: 0 B: 0
		188 =>	x"00000000", -- R: 0 G: 0 B: 0
		189 =>	x"00000000", -- R: 0 G: 0 B: 0
		190 =>	x"00000000", -- R: 0 G: 0 B: 0
		191 =>	x"00000000", -- R: 0 G: 0 B: 0
		192 =>	x"00000000", -- R: 0 G: 0 B: 0
		193 =>	x"00000000", -- R: 0 G: 0 B: 0
		194 =>	x"00000000", -- R: 0 G: 0 B: 0
		195 =>	x"00000000", -- R: 0 G: 0 B: 0
		196 =>	x"00000000", -- R: 0 G: 0 B: 0
		197 =>	x"00000000", -- R: 0 G: 0 B: 0
		198 =>	x"00000000", -- R: 0 G: 0 B: 0
		199 =>	x"00000000", -- R: 0 G: 0 B: 0
		200 =>	x"00000000", -- R: 0 G: 0 B: 0
		201 =>	x"00000000", -- R: 0 G: 0 B: 0
		202 =>	x"00000000", -- R: 0 G: 0 B: 0
		203 =>	x"00000000", -- R: 0 G: 0 B: 0
		204 =>	x"00000000", -- R: 0 G: 0 B: 0
		205 =>	x"00000000", -- R: 0 G: 0 B: 0
		206 =>	x"00000000", -- R: 0 G: 0 B: 0
		207 =>	x"00000000", -- R: 0 G: 0 B: 0
		208 =>	x"00000000", -- R: 0 G: 0 B: 0
		209 =>	x"00000000", -- R: 0 G: 0 B: 0
		210 =>	x"00000000", -- R: 0 G: 0 B: 0
		211 =>	x"00000000", -- R: 0 G: 0 B: 0
		212 =>	x"00000000", -- R: 0 G: 0 B: 0
		213 =>	x"00000000", -- R: 0 G: 0 B: 0
		214 =>	x"00000000", -- R: 0 G: 0 B: 0
		215 =>	x"00000000", -- R: 0 G: 0 B: 0
		216 =>	x"00000000", -- R: 0 G: 0 B: 0
		217 =>	x"00000000", -- R: 0 G: 0 B: 0
		218 =>	x"00000000", -- R: 0 G: 0 B: 0
		219 =>	x"00000000", -- R: 0 G: 0 B: 0
		220 =>	x"00000000", -- R: 0 G: 0 B: 0
		221 =>	x"00000000", -- R: 0 G: 0 B: 0
		222 =>	x"00000000", -- R: 0 G: 0 B: 0
		223 =>	x"00000000", -- R: 0 G: 0 B: 0
		224 =>	x"00000000", -- R: 0 G: 0 B: 0
		225 =>	x"00000000", -- R: 0 G: 0 B: 0
		226 =>	x"00000000", -- R: 0 G: 0 B: 0
		227 =>	x"00000000", -- R: 0 G: 0 B: 0
		228 =>	x"00000000", -- R: 0 G: 0 B: 0
		229 =>	x"00000000", -- R: 0 G: 0 B: 0
		230 =>	x"00000000", -- R: 0 G: 0 B: 0
		231 =>	x"00000000", -- R: 0 G: 0 B: 0
		232 =>	x"00000000", -- R: 0 G: 0 B: 0
		233 =>	x"00000000", -- R: 0 G: 0 B: 0
		234 =>	x"00000000", -- R: 0 G: 0 B: 0
		235 =>	x"00000000", -- R: 0 G: 0 B: 0
		236 =>	x"00000000", -- R: 0 G: 0 B: 0
		237 =>	x"00000000", -- R: 0 G: 0 B: 0
		238 =>	x"00000000", -- R: 0 G: 0 B: 0
		239 =>	x"00000000", -- R: 0 G: 0 B: 0
		240 =>	x"00000000", -- R: 0 G: 0 B: 0
		241 =>	x"00000000", -- R: 0 G: 0 B: 0
		242 =>	x"00000000", -- R: 0 G: 0 B: 0
		243 =>	x"00000000", -- R: 0 G: 0 B: 0
		244 =>	x"00000000", -- R: 0 G: 0 B: 0
		245 =>	x"00000000", -- R: 0 G: 0 B: 0
		246 =>	x"00000000", -- R: 0 G: 0 B: 0
		247 =>	x"00000000", -- R: 0 G: 0 B: 0
		248 =>	x"00000000", -- R: 0 G: 0 B: 0
		249 =>	x"00000000", -- R: 0 G: 0 B: 0
		250 =>	x"00000000", -- R: 0 G: 0 B: 0
		251 =>	x"00000000", -- R: 0 G: 0 B: 0
		252 =>	x"00000000", -- R: 0 G: 0 B: 0
		253 =>	x"00000000", -- R: 0 G: 0 B: 0
		254 =>	x"00000000", -- R: 0 G: 0 B: 0
		255 =>	x"00000000", -- R: 0 G: 0 B: 0


--			***** 16x16 IMAGES *****


		255 =>	x"01020202", -- IMG_16x16_cigle
		256 =>	x"02020202",
		257 =>	x"02000102",
		258 =>	x"02020201",
		259 =>	x"02010101",
		260 =>	x"01010101",
		261 =>	x"01000201",
		262 =>	x"01010100",
		263 =>	x"02010101",
		264 =>	x"01010101",
		265 =>	x"01000201",
		266 =>	x"01010100",
		267 =>	x"02010101",
		268 =>	x"01010101",
		269 =>	x"01000201",
		270 =>	x"01010100",
		271 =>	x"02010101",
		272 =>	x"01010101",
		273 =>	x"01000200",
		274 =>	x"01010100",
		275 =>	x"02010101",
		276 =>	x"01010101",
		277 =>	x"01000100",
		278 =>	x"00000001",
		279 =>	x"02010101",
		280 =>	x"01010101",
		281 =>	x"01000202",
		282 =>	x"02020200",
		283 =>	x"02010101",
		284 =>	x"01010101",
		285 =>	x"01000201",
		286 =>	x"01010100",
		287 =>	x"02010101",
		288 =>	x"01010101",
		289 =>	x"01000201",
		290 =>	x"01010100",
		291 =>	x"02010101",
		292 =>	x"01010101",
		293 =>	x"01000201",
		294 =>	x"01010100",
		295 =>	x"00000101",
		296 =>	x"01010101",
		297 =>	x"00020101",
		298 =>	x"01010100",
		299 =>	x"02020000",
		300 =>	x"01010101",
		301 =>	x"00020101",
		302 =>	x"01010100",
		303 =>	x"02010202",
		304 =>	x"00000000",
		305 =>	x"02010101",
		306 =>	x"01010100",
		307 =>	x"02010101",
		308 =>	x"02020200",
		309 =>	x"02010101",
		310 =>	x"01010100",
		311 =>	x"02010101",
		312 =>	x"01010100",
		313 =>	x"02010101",
		314 =>	x"01010000",
		315 =>	x"01000000",
		316 =>	x"00000001",
		317 =>	x"02000000",
		318 =>	x"00000001",
		319 =>	x"03030304", -- IMG_16x16_coin
		320 =>	x"05060707",
		321 =>	x"08090A0B",
		322 =>	x"0C030303",
		323 =>	x"0303030D",
		324 =>	x"0E0F100F",
		325 =>	x"11121314",
		326 =>	x"15030303",
		327 =>	x"03031617",
		328 =>	x"18191A1B",
		329 =>	x"1C1D1E1F",
		330 =>	x"20210303",
		331 =>	x"22230724",
		332 =>	x"25262728",
		333 =>	x"292A2B2B",
		334 =>	x"2C2D2E2F",
		335 =>	x"30300731",
		336 =>	x"32183033",
		337 =>	x"342D2B35",
		338 =>	x"362D2D2D",
		339 =>	x"30300731",
		340 =>	x"32183033",
		341 =>	x"342D2B35",
		342 =>	x"362D2D2D",
		343 =>	x"30300731",
		344 =>	x"32183033",
		345 =>	x"342D2B35",
		346 =>	x"362D2D2D",
		347 =>	x"30300731",
		348 =>	x"32183033",
		349 =>	x"342D2B35",
		350 =>	x"362D2D2D",
		351 =>	x"30300731",
		352 =>	x"32183033",
		353 =>	x"342D2B35",
		354 =>	x"362D2D2D",
		355 =>	x"30300731",
		356 =>	x"32183033",
		357 =>	x"342D2B35",
		358 =>	x"362D2D2D",
		359 =>	x"30300731",
		360 =>	x"32183033",
		361 =>	x"342D2B35",
		362 =>	x"362D2D2D",
		363 =>	x"30300731",
		364 =>	x"32183033",
		365 =>	x"342D2B35",
		366 =>	x"362D2D2D",
		367 =>	x"22230724",
		368 =>	x"25373338",
		369 =>	x"392A2B2B",
		370 =>	x"2C2D2E2F",
		371 =>	x"03031617",
		372 =>	x"3A0A3B0A",
		373 =>	x"3C3D1E1F",
		374 =>	x"20210303",
		375 =>	x"0303033E",
		376 =>	x"3F404142",
		377 =>	x"43441314",
		378 =>	x"15030303",
		379 =>	x"03030304",
		380 =>	x"05454545",
		381 =>	x"46470A0B",
		382 =>	x"0C030303",
		383 =>	x"48484848", -- IMG_16x16_crno
		384 =>	x"48484848",
		385 =>	x"48484848",
		386 =>	x"48484848",
		387 =>	x"48484848",
		388 =>	x"48484848",
		389 =>	x"48484848",
		390 =>	x"48484848",
		391 =>	x"48484848",
		392 =>	x"48484848",
		393 =>	x"48484848",
		394 =>	x"48484848",
		395 =>	x"48484848",
		396 =>	x"48484848",
		397 =>	x"48484848",
		398 =>	x"48484848",
		399 =>	x"48484848",
		400 =>	x"48484848",
		401 =>	x"48484848",
		402 =>	x"48484848",
		403 =>	x"48484848",
		404 =>	x"48484848",
		405 =>	x"48484848",
		406 =>	x"48484848",
		407 =>	x"48484848",
		408 =>	x"48484848",
		409 =>	x"48484848",
		410 =>	x"48484848",
		411 =>	x"48484848",
		412 =>	x"48484848",
		413 =>	x"48484848",
		414 =>	x"48484848",
		415 =>	x"48484848",
		416 =>	x"48484848",
		417 =>	x"48484848",
		418 =>	x"48484848",
		419 =>	x"48484848",
		420 =>	x"48484848",
		421 =>	x"48484848",
		422 =>	x"48484848",
		423 =>	x"48484848",
		424 =>	x"48484848",
		425 =>	x"48484848",
		426 =>	x"48484848",
		427 =>	x"48484848",
		428 =>	x"48484848",
		429 =>	x"48484848",
		430 =>	x"48484848",
		431 =>	x"48484848",
		432 =>	x"48484848",
		433 =>	x"48484848",
		434 =>	x"48484848",
		435 =>	x"48484848",
		436 =>	x"48484848",
		437 =>	x"48484848",
		438 =>	x"48484848",
		439 =>	x"48484848",
		440 =>	x"48484848",
		441 =>	x"48484848",
		442 =>	x"48484848",
		443 =>	x"48484848",
		444 =>	x"48484848",
		445 =>	x"48484848",
		446 =>	x"48484848",
		447 =>	x"03030303", -- IMG_16x16_enemi1
		448 =>	x"03494949",
		449 =>	x"49490303",
		450 =>	x"03030303",
		451 =>	x"03030303",
		452 =>	x"49494949",
		453 =>	x"49494903",
		454 =>	x"03030303",
		455 =>	x"03030349",
		456 =>	x"49494949",
		457 =>	x"49494949",
		458 =>	x"03030303",
		459 =>	x"03034949",
		460 =>	x"49494949",
		461 =>	x"49494949",
		462 =>	x"49030303",
		463 =>	x"03494A4A",
		464 =>	x"49494949",
		465 =>	x"4949494A",
		466 =>	x"4A490303",
		467 =>	x"4949494B",
		468 =>	x"4A494949",
		469 =>	x"49494A4B",
		470 =>	x"49494903",
		471 =>	x"4949494B",
		472 =>	x"4A4A4A4A",
		473 =>	x"4A4A4A4B",
		474 =>	x"49494903",
		475 =>	x"4949494B",
		476 =>	x"4A4B4949",
		477 =>	x"494B4A4B",
		478 =>	x"49494949",
		479 =>	x"4949494B",
		480 =>	x"4B4B4949",
		481 =>	x"494B4B4B",
		482 =>	x"49494949",
		483 =>	x"49494949",
		484 =>	x"49494949",
		485 =>	x"49494949",
		486 =>	x"49494949",
		487 =>	x"49494949",
		488 =>	x"4B4B4B4B",
		489 =>	x"4B4B4B49",
		490 =>	x"49494903",
		491 =>	x"0303034B",
		492 =>	x"4B4B4B4B",
		493 =>	x"4B4B4B4B",
		494 =>	x"03030303",
		495 =>	x"0300004B",
		496 =>	x"4B4B4B4B",
		497 =>	x"4B4B4B4B",
		498 =>	x"03030303",
		499 =>	x"00000000",
		500 =>	x"004B4B4B",
		501 =>	x"4B4B4B00",
		502 =>	x"00030303",
		503 =>	x"00000000",
		504 =>	x"00004B4B",
		505 =>	x"4B4B0000",
		506 =>	x"00030303",
		507 =>	x"03000000",
		508 =>	x"00000303",
		509 =>	x"03000000",
		510 =>	x"03030303",
		511 =>	x"03034C4C", -- IMG_16x16_mario
		512 =>	x"4C4C4C4C",
		513 =>	x"4C4C4C4C",
		514 =>	x"4C4C4C03",
		515 =>	x"03034D4D",
		516 =>	x"4D4D4E4E",
		517 =>	x"4E4D4E4E",
		518 =>	x"03030303",
		519 =>	x"034D4E4E",
		520 =>	x"4D4E4E4E",
		521 =>	x"4E4D4F4E",
		522 =>	x"4E4E4E03",
		523 =>	x"034D5050",
		524 =>	x"4D4D4E4E",
		525 =>	x"4E4F4D4E",
		526 =>	x"4E4E4E4E",
		527 =>	x"034D4D4D",
		528 =>	x"514E4E4E",
		529 =>	x"4E4D4D4D",
		530 =>	x"4D4D4D03",
		531 =>	x"03030303",
		532 =>	x"4E4E4E4E",
		533 =>	x"4E4E4E4E",
		534 =>	x"4E4E0303",
		535 =>	x"03034D4D",
		536 =>	x"4D4C4D4D",
		537 =>	x"4D4D4D03",
		538 =>	x"03030303",
		539 =>	x"034D4D4D",
		540 =>	x"4D4C4D4D",
		541 =>	x"4D4C4D4D",
		542 =>	x"4D4D4D03",
		543 =>	x"034D4D4D",
		544 =>	x"4D4C4D4D",
		545 =>	x"4D4C4D4D",
		546 =>	x"4D4D4D03",
		547 =>	x"4D4D4D4D",
		548 =>	x"4D4C4C4C",
		549 =>	x"4C4C4D4D",
		550 =>	x"4D4D4D4D",
		551 =>	x"4E4E4D4D",
		552 =>	x"4C4E4C4C",
		553 =>	x"4C4E4C4D",
		554 =>	x"4E4E4E4E",
		555 =>	x"4E4E4E4E",
		556 =>	x"4C4C4C4C",
		557 =>	x"4C4C4C4E",
		558 =>	x"4E4E4E4E",
		559 =>	x"4E4E4C4C",
		560 =>	x"4C4C4C4C",
		561 =>	x"4C4C4C4C",
		562 =>	x"4E4E4E4E",
		563 =>	x"03034C4C",
		564 =>	x"4C4C4C03",
		565 =>	x"034C4C4C",
		566 =>	x"4C4C0303",
		567 =>	x"034D4D4D",
		568 =>	x"4D4D0303",
		569 =>	x"03034D4D",
		570 =>	x"4D4D4D03",
		571 =>	x"4D4D4D4D",
		572 =>	x"4D4D0303",
		573 =>	x"03034D4D",
		574 =>	x"4D4D4D4D",
		575 =>	x"00000000", -- IMG_16x16_plavacigla
		576 =>	x"00000000",
		577 =>	x"00000000",
		578 =>	x"00000000",
		579 =>	x"49494949",
		580 =>	x"49494900",
		581 =>	x"49494949",
		582 =>	x"49494900",
		583 =>	x"49494949",
		584 =>	x"49494900",
		585 =>	x"49494949",
		586 =>	x"49494900",
		587 =>	x"00000000",
		588 =>	x"00000000",
		589 =>	x"00000000",
		590 =>	x"00000000",
		591 =>	x"49494900",
		592 =>	x"49494949",
		593 =>	x"49494900",
		594 =>	x"49494949",
		595 =>	x"49494900",
		596 =>	x"49494949",
		597 =>	x"49494900",
		598 =>	x"49494949",
		599 =>	x"49494900",
		600 =>	x"49494949",
		601 =>	x"49494900",
		602 =>	x"49494949",
		603 =>	x"00000000",
		604 =>	x"00000000",
		605 =>	x"00000000",
		606 =>	x"00000000",
		607 =>	x"49494949",
		608 =>	x"49494900",
		609 =>	x"49494949",
		610 =>	x"49494900",
		611 =>	x"49494949",
		612 =>	x"49494900",
		613 =>	x"49494949",
		614 =>	x"49494900",
		615 =>	x"49494949",
		616 =>	x"49494900",
		617 =>	x"49494949",
		618 =>	x"49494900",
		619 =>	x"00000000",
		620 =>	x"00000000",
		621 =>	x"00000000",
		622 =>	x"00000000",
		623 =>	x"49494900",
		624 =>	x"49494949",
		625 =>	x"49494900",
		626 =>	x"49494949",
		627 =>	x"49494900",
		628 =>	x"49494949",
		629 =>	x"49494900",
		630 =>	x"49494949",
		631 =>	x"49494900",
		632 =>	x"49494949",
		633 =>	x"49494900",
		634 =>	x"49494949",
		635 =>	x"00000000",
		636 =>	x"00000000",
		637 =>	x"00000000",
		638 =>	x"00000000",


--			***** MAP *****


		639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		1999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2879 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2880 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2881 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2882 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2883 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2884 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2885 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2886 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2887 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2888 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2889 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2890 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2891 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2892 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2893 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2894 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2895 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2896 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2897 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2898 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2899 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2900 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2901 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2902 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2903 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2904 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2905 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2906 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2907 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2908 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2909 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2910 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2911 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2912 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2913 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2914 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2915 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2916 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2917 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2918 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2919 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2959 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2960 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2961 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2962 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2963 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2964 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2965 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2966 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2967 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2968 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2969 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2970 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2971 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2972 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2973 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2974 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2975 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2976 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2977 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2978 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2979 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2980 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2981 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2982 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2983 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2984 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2985 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2986 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2987 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2988 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2989 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2990 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2991 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2992 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2993 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2994 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2995 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2996 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2997 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2998 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		2999 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		3000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3199 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3583 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"
	);



		
begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;